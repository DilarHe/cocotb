// Generator : SpinalHDL v1.8.0    git head : 4e3563a282582b41f4eaafc503787757251d23ea
// Component : registers
// Git hash  : a8f29ef6fd0b904c29693408b375c85f91553a49

`timescale 1ns/1ps 
module registers (
  input      [4:0]    dec_rs1_index,
  input      [4:0]    dec_rs2_index,
  input      [4:0]    dec_rd_index,
  input      [31:0]   dec_imm,
  input               dec_imm_is_rs2,
  input               dec_is_jump,
  input               dec_is_branch,
  input               dec_is_wload,
  input               dec_is_wstore,
  input               dec_is_multi_rs1_index,
  input               dec_is_vector_oprand_used,
  input               dec_is_vload,
  input               dec_is_vstore1,
  input               dec_is_vstore2,
  input               dec_info_vld,
  input      [31:0]   alu_write_rd_data,
  input      [4:0]    alu_write_rd_index,
  input               alu_write_rd_vld,
  input      [31:0]   lsu_write_rd_data,
  input      [4:0]    lsu_write_rd_index,
  input               lsu_write_rd_vld,
  input               lsu_write_rd_is_vector,
  input      [127:0]  lsu_write_rd_vector_data,
  output     [31:0]   roperand_out_rs1,
  output     [4:0]    roperand_out_rs1_index,
  output     [31:0]   roperand_out_rs2,
  output     [4:0]    roperand_out_rs2_index,
  output     [4:0]    roperand_out_rd_index,
  output reg [127:0]  voperand_out_vs1,
  output reg [127:0]  voperand_out_vs2,
  output     [4:0]    voperand_out_vs1_index,
  output     [4:0]    voperand_out_vs2_index,
  output              oprand_vld_out,
  input               clk,
  input               resetn
);

  reg        [31:0]   tmp_tmp_roperand_out_rs1;
  reg        [31:0]   tmp_roperand_out_rs1_1;
  wire       [4:0]    tmp_roperand_out_rs1_2;
  reg        [31:0]   tmp_roperand_out_rs2;
  reg        [31:0]   tmp_roperand_out_rd_index;
  wire                lsu_write_normal_regfile_vld;
  wire                lsu_write_vector_regfile_vld;
  wire       [4:0]    lsu_write_normal_rd_index;
  wire       [31:0]   lsu_write_normal_rd_data;
  wire       [4:0]    write_vector_rd_index_0;
  wire       [4:0]    write_vector_rd_index_1;
  wire       [4:0]    write_vector_rd_index_2;
  wire       [4:0]    write_vector_rd_index_3;
  wire       [31:0]   write_vector_rd_data_0;
  wire       [31:0]   write_vector_rd_data_1;
  wire       [31:0]   write_vector_rd_data_2;
  wire       [31:0]   write_vector_rd_data_3;
  reg        [31:0]   x_0;
  reg        [31:0]   x_1;
  reg        [31:0]   x_2;
  reg        [31:0]   x_3;
  reg        [31:0]   x_4;
  reg        [31:0]   x_5;
  reg        [31:0]   x_6;
  reg        [31:0]   x_7;
  reg        [31:0]   x_8;
  reg        [31:0]   x_9;
  reg        [31:0]   x_10;
  reg        [31:0]   x_11;
  reg        [31:0]   x_12;
  reg        [31:0]   x_13;
  reg        [31:0]   x_14;
  reg        [31:0]   x_15;
  reg        [31:0]   x_16;
  reg        [31:0]   x_17;
  reg        [31:0]   x_18;
  reg        [31:0]   x_19;
  reg        [31:0]   x_20;
  reg        [31:0]   x_21;
  reg        [31:0]   x_22;
  reg        [31:0]   x_23;
  reg        [31:0]   x_24;
  reg        [31:0]   x_25;
  reg        [31:0]   x_26;
  reg        [31:0]   x_27;
  reg        [31:0]   x_28;
  reg        [31:0]   x_29;
  reg        [31:0]   x_30;
  reg        [31:0]   x_31;
  wire       [4:0]    vs2_index;
  wire       [31:0]   tmp_roperand_out_rs1;
  wire                is_vector_instr;

  assign tmp_roperand_out_rs1_2 = tmp_roperand_out_rs1[4 : 0];
  always @(*) begin
    case(dec_rs1_index)
      5'b00000 : tmp_tmp_roperand_out_rs1 = x_0;
      5'b00001 : tmp_tmp_roperand_out_rs1 = x_1;
      5'b00010 : tmp_tmp_roperand_out_rs1 = x_2;
      5'b00011 : tmp_tmp_roperand_out_rs1 = x_3;
      5'b00100 : tmp_tmp_roperand_out_rs1 = x_4;
      5'b00101 : tmp_tmp_roperand_out_rs1 = x_5;
      5'b00110 : tmp_tmp_roperand_out_rs1 = x_6;
      5'b00111 : tmp_tmp_roperand_out_rs1 = x_7;
      5'b01000 : tmp_tmp_roperand_out_rs1 = x_8;
      5'b01001 : tmp_tmp_roperand_out_rs1 = x_9;
      5'b01010 : tmp_tmp_roperand_out_rs1 = x_10;
      5'b01011 : tmp_tmp_roperand_out_rs1 = x_11;
      5'b01100 : tmp_tmp_roperand_out_rs1 = x_12;
      5'b01101 : tmp_tmp_roperand_out_rs1 = x_13;
      5'b01110 : tmp_tmp_roperand_out_rs1 = x_14;
      5'b01111 : tmp_tmp_roperand_out_rs1 = x_15;
      5'b10000 : tmp_tmp_roperand_out_rs1 = x_16;
      5'b10001 : tmp_tmp_roperand_out_rs1 = x_17;
      5'b10010 : tmp_tmp_roperand_out_rs1 = x_18;
      5'b10011 : tmp_tmp_roperand_out_rs1 = x_19;
      5'b10100 : tmp_tmp_roperand_out_rs1 = x_20;
      5'b10101 : tmp_tmp_roperand_out_rs1 = x_21;
      5'b10110 : tmp_tmp_roperand_out_rs1 = x_22;
      5'b10111 : tmp_tmp_roperand_out_rs1 = x_23;
      5'b11000 : tmp_tmp_roperand_out_rs1 = x_24;
      5'b11001 : tmp_tmp_roperand_out_rs1 = x_25;
      5'b11010 : tmp_tmp_roperand_out_rs1 = x_26;
      5'b11011 : tmp_tmp_roperand_out_rs1 = x_27;
      5'b11100 : tmp_tmp_roperand_out_rs1 = x_28;
      5'b11101 : tmp_tmp_roperand_out_rs1 = x_29;
      5'b11110 : tmp_tmp_roperand_out_rs1 = x_30;
      default : tmp_tmp_roperand_out_rs1 = x_31;
    endcase
  end

  always @(*) begin
    case(tmp_roperand_out_rs1_2)
      5'b00000 : tmp_roperand_out_rs1_1 = x_0;
      5'b00001 : tmp_roperand_out_rs1_1 = x_1;
      5'b00010 : tmp_roperand_out_rs1_1 = x_2;
      5'b00011 : tmp_roperand_out_rs1_1 = x_3;
      5'b00100 : tmp_roperand_out_rs1_1 = x_4;
      5'b00101 : tmp_roperand_out_rs1_1 = x_5;
      5'b00110 : tmp_roperand_out_rs1_1 = x_6;
      5'b00111 : tmp_roperand_out_rs1_1 = x_7;
      5'b01000 : tmp_roperand_out_rs1_1 = x_8;
      5'b01001 : tmp_roperand_out_rs1_1 = x_9;
      5'b01010 : tmp_roperand_out_rs1_1 = x_10;
      5'b01011 : tmp_roperand_out_rs1_1 = x_11;
      5'b01100 : tmp_roperand_out_rs1_1 = x_12;
      5'b01101 : tmp_roperand_out_rs1_1 = x_13;
      5'b01110 : tmp_roperand_out_rs1_1 = x_14;
      5'b01111 : tmp_roperand_out_rs1_1 = x_15;
      5'b10000 : tmp_roperand_out_rs1_1 = x_16;
      5'b10001 : tmp_roperand_out_rs1_1 = x_17;
      5'b10010 : tmp_roperand_out_rs1_1 = x_18;
      5'b10011 : tmp_roperand_out_rs1_1 = x_19;
      5'b10100 : tmp_roperand_out_rs1_1 = x_20;
      5'b10101 : tmp_roperand_out_rs1_1 = x_21;
      5'b10110 : tmp_roperand_out_rs1_1 = x_22;
      5'b10111 : tmp_roperand_out_rs1_1 = x_23;
      5'b11000 : tmp_roperand_out_rs1_1 = x_24;
      5'b11001 : tmp_roperand_out_rs1_1 = x_25;
      5'b11010 : tmp_roperand_out_rs1_1 = x_26;
      5'b11011 : tmp_roperand_out_rs1_1 = x_27;
      5'b11100 : tmp_roperand_out_rs1_1 = x_28;
      5'b11101 : tmp_roperand_out_rs1_1 = x_29;
      5'b11110 : tmp_roperand_out_rs1_1 = x_30;
      default : tmp_roperand_out_rs1_1 = x_31;
    endcase
  end

  always @(*) begin
    case(dec_rs2_index)
      5'b00000 : tmp_roperand_out_rs2 = x_0;
      5'b00001 : tmp_roperand_out_rs2 = x_1;
      5'b00010 : tmp_roperand_out_rs2 = x_2;
      5'b00011 : tmp_roperand_out_rs2 = x_3;
      5'b00100 : tmp_roperand_out_rs2 = x_4;
      5'b00101 : tmp_roperand_out_rs2 = x_5;
      5'b00110 : tmp_roperand_out_rs2 = x_6;
      5'b00111 : tmp_roperand_out_rs2 = x_7;
      5'b01000 : tmp_roperand_out_rs2 = x_8;
      5'b01001 : tmp_roperand_out_rs2 = x_9;
      5'b01010 : tmp_roperand_out_rs2 = x_10;
      5'b01011 : tmp_roperand_out_rs2 = x_11;
      5'b01100 : tmp_roperand_out_rs2 = x_12;
      5'b01101 : tmp_roperand_out_rs2 = x_13;
      5'b01110 : tmp_roperand_out_rs2 = x_14;
      5'b01111 : tmp_roperand_out_rs2 = x_15;
      5'b10000 : tmp_roperand_out_rs2 = x_16;
      5'b10001 : tmp_roperand_out_rs2 = x_17;
      5'b10010 : tmp_roperand_out_rs2 = x_18;
      5'b10011 : tmp_roperand_out_rs2 = x_19;
      5'b10100 : tmp_roperand_out_rs2 = x_20;
      5'b10101 : tmp_roperand_out_rs2 = x_21;
      5'b10110 : tmp_roperand_out_rs2 = x_22;
      5'b10111 : tmp_roperand_out_rs2 = x_23;
      5'b11000 : tmp_roperand_out_rs2 = x_24;
      5'b11001 : tmp_roperand_out_rs2 = x_25;
      5'b11010 : tmp_roperand_out_rs2 = x_26;
      5'b11011 : tmp_roperand_out_rs2 = x_27;
      5'b11100 : tmp_roperand_out_rs2 = x_28;
      5'b11101 : tmp_roperand_out_rs2 = x_29;
      5'b11110 : tmp_roperand_out_rs2 = x_30;
      default : tmp_roperand_out_rs2 = x_31;
    endcase
  end

  always @(*) begin
    case(dec_rd_index)
      5'b00000 : tmp_roperand_out_rd_index = x_0;
      5'b00001 : tmp_roperand_out_rd_index = x_1;
      5'b00010 : tmp_roperand_out_rd_index = x_2;
      5'b00011 : tmp_roperand_out_rd_index = x_3;
      5'b00100 : tmp_roperand_out_rd_index = x_4;
      5'b00101 : tmp_roperand_out_rd_index = x_5;
      5'b00110 : tmp_roperand_out_rd_index = x_6;
      5'b00111 : tmp_roperand_out_rd_index = x_7;
      5'b01000 : tmp_roperand_out_rd_index = x_8;
      5'b01001 : tmp_roperand_out_rd_index = x_9;
      5'b01010 : tmp_roperand_out_rd_index = x_10;
      5'b01011 : tmp_roperand_out_rd_index = x_11;
      5'b01100 : tmp_roperand_out_rd_index = x_12;
      5'b01101 : tmp_roperand_out_rd_index = x_13;
      5'b01110 : tmp_roperand_out_rd_index = x_14;
      5'b01111 : tmp_roperand_out_rd_index = x_15;
      5'b10000 : tmp_roperand_out_rd_index = x_16;
      5'b10001 : tmp_roperand_out_rd_index = x_17;
      5'b10010 : tmp_roperand_out_rd_index = x_18;
      5'b10011 : tmp_roperand_out_rd_index = x_19;
      5'b10100 : tmp_roperand_out_rd_index = x_20;
      5'b10101 : tmp_roperand_out_rd_index = x_21;
      5'b10110 : tmp_roperand_out_rd_index = x_22;
      5'b10111 : tmp_roperand_out_rd_index = x_23;
      5'b11000 : tmp_roperand_out_rd_index = x_24;
      5'b11001 : tmp_roperand_out_rd_index = x_25;
      5'b11010 : tmp_roperand_out_rd_index = x_26;
      5'b11011 : tmp_roperand_out_rd_index = x_27;
      5'b11100 : tmp_roperand_out_rd_index = x_28;
      5'b11101 : tmp_roperand_out_rd_index = x_29;
      5'b11110 : tmp_roperand_out_rd_index = x_30;
      default : tmp_roperand_out_rd_index = x_31;
    endcase
  end

  assign lsu_write_normal_regfile_vld = (lsu_write_rd_vld && (! lsu_write_rd_is_vector)); // @[BaseType.scala 305:24]
  assign lsu_write_vector_regfile_vld = (lsu_write_rd_vld && lsu_write_rd_is_vector); // @[BaseType.scala 305:24]
  assign lsu_write_normal_rd_index = (lsu_write_normal_regfile_vld ? lsu_write_rd_index : 5'h0); // @[Expression.scala 1420:25]
  assign lsu_write_normal_rd_data = (lsu_write_normal_regfile_vld ? lsu_write_rd_data : 32'h0); // @[Expression.scala 1420:25]
  assign write_vector_rd_index_0 = (lsu_write_rd_index + 5'h0); // @[registers.scala 49:30]
  assign write_vector_rd_data_0 = lsu_write_rd_vector_data[31 : 0]; // @[registers.scala 50:29]
  assign write_vector_rd_index_1 = (lsu_write_rd_index + 5'h01); // @[registers.scala 49:30]
  assign write_vector_rd_data_1 = lsu_write_rd_vector_data[63 : 32]; // @[registers.scala 50:29]
  assign write_vector_rd_index_2 = (lsu_write_rd_index + 5'h02); // @[registers.scala 49:30]
  assign write_vector_rd_data_2 = lsu_write_rd_vector_data[95 : 64]; // @[registers.scala 50:29]
  assign write_vector_rd_index_3 = (lsu_write_rd_index + 5'h03); // @[registers.scala 49:30]
  assign write_vector_rd_data_3 = lsu_write_rd_vector_data[127 : 96]; // @[registers.scala 50:29]
  assign vs2_index = (dec_rs2_index + 5'h04); // @[BaseType.scala 299:24]
  assign voperand_out_vs1_index = dec_rs2_index; // @[registers.scala 106:29]
  assign voperand_out_vs2_index = vs2_index; // @[registers.scala 107:29]
  assign tmp_roperand_out_rs1 = tmp_tmp_roperand_out_rs1; // @[Vec.scala 202:25]
  assign roperand_out_rs1_index = (dec_is_multi_rs1_index ? tmp_roperand_out_rs1[4 : 0] : dec_rs1_index); // @[registers.scala 109:29]
  assign roperand_out_rs2_index = (dec_imm_is_rs2 ? 5'h0 : dec_rs2_index); // @[registers.scala 110:29]
  assign roperand_out_rs1 = (dec_is_multi_rs1_index ? tmp_roperand_out_rs1_1 : tmp_roperand_out_rs1); // @[registers.scala 111:23]
  assign roperand_out_rs2 = (dec_imm_is_rs2 ? dec_imm : tmp_roperand_out_rs2); // @[registers.scala 112:23]
  assign roperand_out_rd_index = (dec_is_multi_rs1_index ? tmp_roperand_out_rd_index[4 : 0] : dec_rd_index); // @[registers.scala 113:28]
  assign oprand_vld_out = dec_info_vld; // @[registers.scala 120:21]
  assign is_vector_instr = (((dec_is_vector_oprand_used || dec_is_vload) || dec_is_vstore1) || dec_is_vstore2); // @[BaseType.scala 305:24]
  always @(*) begin
    if(is_vector_instr) begin
      voperand_out_vs1[31 : 0] = x_8; // @[registers.scala 128:59]
      voperand_out_vs1[63 : 32] = x_9; // @[registers.scala 128:59]
      voperand_out_vs1[95 : 64] = x_10; // @[registers.scala 128:59]
      voperand_out_vs1[127 : 96] = x_11; // @[registers.scala 128:59]
    end else begin
      voperand_out_vs1 = 128'h0; // @[registers.scala 131:25]
    end
  end

  always @(*) begin
    if(is_vector_instr) begin
      voperand_out_vs2[31 : 0] = x_12; // @[registers.scala 139:59]
      voperand_out_vs2[63 : 32] = x_13; // @[registers.scala 139:59]
      voperand_out_vs2[95 : 64] = x_14; // @[registers.scala 139:59]
      voperand_out_vs2[127 : 96] = x_15; // @[registers.scala 139:59]
    end else begin
      if(dec_is_vstore1) begin
        voperand_out_vs2[7 : 0] = x_16[7 : 0]; // @[registers.scala 143:73]
        voperand_out_vs2[15 : 8] = x_17[7 : 0]; // @[registers.scala 143:73]
        voperand_out_vs2[23 : 16] = x_18[7 : 0]; // @[registers.scala 143:73]
        voperand_out_vs2[31 : 24] = x_19[7 : 0]; // @[registers.scala 143:73]
        voperand_out_vs2[39 : 32] = x_20[7 : 0]; // @[registers.scala 143:73]
        voperand_out_vs2[47 : 40] = x_21[7 : 0]; // @[registers.scala 143:73]
        voperand_out_vs2[55 : 48] = x_22[7 : 0]; // @[registers.scala 143:73]
        voperand_out_vs2[63 : 56] = x_23[7 : 0]; // @[registers.scala 143:73]
        voperand_out_vs2[71 : 64] = x_24[7 : 0]; // @[registers.scala 143:73]
        voperand_out_vs2[79 : 72] = x_25[7 : 0]; // @[registers.scala 143:73]
        voperand_out_vs2[87 : 80] = x_26[7 : 0]; // @[registers.scala 143:73]
        voperand_out_vs2[95 : 88] = x_27[7 : 0]; // @[registers.scala 143:73]
        voperand_out_vs2[103 : 96] = x_28[7 : 0]; // @[registers.scala 143:73]
        voperand_out_vs2[111 : 104] = x_29[7 : 0]; // @[registers.scala 143:73]
        voperand_out_vs2[119 : 112] = x_30[7 : 0]; // @[registers.scala 143:73]
        voperand_out_vs2[127 : 120] = x_31[7 : 0]; // @[registers.scala 143:73]
      end else begin
        voperand_out_vs2 = 128'h0; // @[registers.scala 152:25]
      end
    end
  end

  always @(posedge clk or negedge resetn) begin
    if(!resetn) begin
      x_0 <= 32'h0; // @[Data.scala 400:33]
      x_1 <= 32'h0; // @[Data.scala 400:33]
      x_2 <= 32'h0; // @[Data.scala 400:33]
      x_3 <= 32'h0; // @[Data.scala 400:33]
      x_4 <= 32'h0; // @[Data.scala 400:33]
      x_5 <= 32'h0; // @[Data.scala 400:33]
      x_6 <= 32'h0; // @[Data.scala 400:33]
      x_7 <= 32'h0; // @[Data.scala 400:33]
      x_8 <= 32'h0; // @[Data.scala 400:33]
      x_9 <= 32'h0; // @[Data.scala 400:33]
      x_10 <= 32'h0; // @[Data.scala 400:33]
      x_11 <= 32'h0; // @[Data.scala 400:33]
      x_12 <= 32'h0; // @[Data.scala 400:33]
      x_13 <= 32'h0; // @[Data.scala 400:33]
      x_14 <= 32'h0; // @[Data.scala 400:33]
      x_15 <= 32'h0; // @[Data.scala 400:33]
      x_16 <= 32'h0; // @[Data.scala 400:33]
      x_17 <= 32'h0; // @[Data.scala 400:33]
      x_18 <= 32'h0; // @[Data.scala 400:33]
      x_19 <= 32'h0; // @[Data.scala 400:33]
      x_20 <= 32'h0; // @[Data.scala 400:33]
      x_21 <= 32'h0; // @[Data.scala 400:33]
      x_22 <= 32'h0; // @[Data.scala 400:33]
      x_23 <= 32'h0; // @[Data.scala 400:33]
      x_24 <= 32'h0; // @[Data.scala 400:33]
      x_25 <= 32'h0; // @[Data.scala 400:33]
      x_26 <= 32'h0; // @[Data.scala 400:33]
      x_27 <= 32'h0; // @[Data.scala 400:33]
      x_28 <= 32'h0; // @[Data.scala 400:33]
      x_29 <= 32'h0; // @[Data.scala 400:33]
      x_30 <= 32'h0; // @[Data.scala 400:33]
      x_31 <= 32'h0; // @[Data.scala 400:33]
    end else begin
      x_0 <= 32'h0; // @[registers.scala 55:8]
      if((alu_write_rd_vld && (alu_write_rd_index == 5'h01))) begin
        x_1 <= alu_write_rd_data; // @[registers.scala 72:14]
      end else begin
        if((lsu_write_normal_regfile_vld && (lsu_write_normal_rd_index == 5'h01))) begin
          x_1 <= lsu_write_normal_rd_data; // @[registers.scala 74:14]
        end
      end
      if((alu_write_rd_vld && (alu_write_rd_index == 5'h02))) begin
        x_2 <= alu_write_rd_data; // @[registers.scala 72:14]
      end else begin
        if((lsu_write_normal_regfile_vld && (lsu_write_normal_rd_index == 5'h02))) begin
          x_2 <= lsu_write_normal_rd_data; // @[registers.scala 74:14]
        end
      end
      if((alu_write_rd_vld && (alu_write_rd_index == 5'h03))) begin
        x_3 <= alu_write_rd_data; // @[registers.scala 72:14]
      end else begin
        if((lsu_write_normal_regfile_vld && (lsu_write_normal_rd_index == 5'h03))) begin
          x_3 <= lsu_write_normal_rd_data; // @[registers.scala 74:14]
        end
      end
      if((alu_write_rd_vld && (alu_write_rd_index == 5'h04))) begin
        x_4 <= alu_write_rd_data; // @[registers.scala 72:14]
      end else begin
        if((lsu_write_normal_regfile_vld && (lsu_write_normal_rd_index == 5'h04))) begin
          x_4 <= lsu_write_normal_rd_data; // @[registers.scala 74:14]
        end
      end
      if((alu_write_rd_vld && (alu_write_rd_index == 5'h05))) begin
        x_5 <= alu_write_rd_data; // @[registers.scala 72:14]
      end else begin
        if((lsu_write_normal_regfile_vld && (lsu_write_normal_rd_index == 5'h05))) begin
          x_5 <= lsu_write_normal_rd_data; // @[registers.scala 74:14]
        end
      end
      if((alu_write_rd_vld && (alu_write_rd_index == 5'h06))) begin
        x_6 <= alu_write_rd_data; // @[registers.scala 72:14]
      end else begin
        if((lsu_write_normal_regfile_vld && (lsu_write_normal_rd_index == 5'h06))) begin
          x_6 <= lsu_write_normal_rd_data; // @[registers.scala 74:14]
        end
      end
      if((alu_write_rd_vld && (alu_write_rd_index == 5'h07))) begin
        x_7 <= alu_write_rd_data; // @[registers.scala 72:14]
      end else begin
        if((lsu_write_normal_regfile_vld && (lsu_write_normal_rd_index == 5'h07))) begin
          x_7 <= lsu_write_normal_rd_data; // @[registers.scala 74:14]
        end
      end
      if((alu_write_rd_vld && (alu_write_rd_index == 5'h08))) begin
        x_8 <= alu_write_rd_data; // @[registers.scala 79:14]
      end else begin
        if((lsu_write_normal_regfile_vld && (lsu_write_normal_rd_index == 5'h08))) begin
          x_8 <= lsu_write_normal_rd_data; // @[registers.scala 81:14]
        end else begin
          if(lsu_write_vector_regfile_vld) begin
            if((write_vector_rd_index_0 == 5'h08)) begin
              x_8 <= write_vector_rd_data_0; // @[registers.scala 85:18]
            end
            if((write_vector_rd_index_1 == 5'h08)) begin
              x_8 <= write_vector_rd_data_1; // @[registers.scala 85:18]
            end
            if((write_vector_rd_index_2 == 5'h08)) begin
              x_8 <= write_vector_rd_data_2; // @[registers.scala 85:18]
            end
            if((write_vector_rd_index_3 == 5'h08)) begin
              x_8 <= write_vector_rd_data_3; // @[registers.scala 85:18]
            end
          end
        end
      end
      if((alu_write_rd_vld && (alu_write_rd_index == 5'h09))) begin
        x_9 <= alu_write_rd_data; // @[registers.scala 79:14]
      end else begin
        if((lsu_write_normal_regfile_vld && (lsu_write_normal_rd_index == 5'h09))) begin
          x_9 <= lsu_write_normal_rd_data; // @[registers.scala 81:14]
        end else begin
          if(lsu_write_vector_regfile_vld) begin
            if((write_vector_rd_index_0 == 5'h09)) begin
              x_9 <= write_vector_rd_data_0; // @[registers.scala 85:18]
            end
            if((write_vector_rd_index_1 == 5'h09)) begin
              x_9 <= write_vector_rd_data_1; // @[registers.scala 85:18]
            end
            if((write_vector_rd_index_2 == 5'h09)) begin
              x_9 <= write_vector_rd_data_2; // @[registers.scala 85:18]
            end
            if((write_vector_rd_index_3 == 5'h09)) begin
              x_9 <= write_vector_rd_data_3; // @[registers.scala 85:18]
            end
          end
        end
      end
      if((alu_write_rd_vld && (alu_write_rd_index == 5'h0a))) begin
        x_10 <= alu_write_rd_data; // @[registers.scala 79:14]
      end else begin
        if((lsu_write_normal_regfile_vld && (lsu_write_normal_rd_index == 5'h0a))) begin
          x_10 <= lsu_write_normal_rd_data; // @[registers.scala 81:14]
        end else begin
          if(lsu_write_vector_regfile_vld) begin
            if((write_vector_rd_index_0 == 5'h0a)) begin
              x_10 <= write_vector_rd_data_0; // @[registers.scala 85:18]
            end
            if((write_vector_rd_index_1 == 5'h0a)) begin
              x_10 <= write_vector_rd_data_1; // @[registers.scala 85:18]
            end
            if((write_vector_rd_index_2 == 5'h0a)) begin
              x_10 <= write_vector_rd_data_2; // @[registers.scala 85:18]
            end
            if((write_vector_rd_index_3 == 5'h0a)) begin
              x_10 <= write_vector_rd_data_3; // @[registers.scala 85:18]
            end
          end
        end
      end
      if((alu_write_rd_vld && (alu_write_rd_index == 5'h0b))) begin
        x_11 <= alu_write_rd_data; // @[registers.scala 79:14]
      end else begin
        if((lsu_write_normal_regfile_vld && (lsu_write_normal_rd_index == 5'h0b))) begin
          x_11 <= lsu_write_normal_rd_data; // @[registers.scala 81:14]
        end else begin
          if(lsu_write_vector_regfile_vld) begin
            if((write_vector_rd_index_0 == 5'h0b)) begin
              x_11 <= write_vector_rd_data_0; // @[registers.scala 85:18]
            end
            if((write_vector_rd_index_1 == 5'h0b)) begin
              x_11 <= write_vector_rd_data_1; // @[registers.scala 85:18]
            end
            if((write_vector_rd_index_2 == 5'h0b)) begin
              x_11 <= write_vector_rd_data_2; // @[registers.scala 85:18]
            end
            if((write_vector_rd_index_3 == 5'h0b)) begin
              x_11 <= write_vector_rd_data_3; // @[registers.scala 85:18]
            end
          end
        end
      end
      if((alu_write_rd_vld && (alu_write_rd_index == 5'h0c))) begin
        x_12 <= alu_write_rd_data; // @[registers.scala 79:14]
      end else begin
        if((lsu_write_normal_regfile_vld && (lsu_write_normal_rd_index == 5'h0c))) begin
          x_12 <= lsu_write_normal_rd_data; // @[registers.scala 81:14]
        end else begin
          if(lsu_write_vector_regfile_vld) begin
            if((write_vector_rd_index_0 == 5'h0c)) begin
              x_12 <= write_vector_rd_data_0; // @[registers.scala 85:18]
            end
            if((write_vector_rd_index_1 == 5'h0c)) begin
              x_12 <= write_vector_rd_data_1; // @[registers.scala 85:18]
            end
            if((write_vector_rd_index_2 == 5'h0c)) begin
              x_12 <= write_vector_rd_data_2; // @[registers.scala 85:18]
            end
            if((write_vector_rd_index_3 == 5'h0c)) begin
              x_12 <= write_vector_rd_data_3; // @[registers.scala 85:18]
            end
          end
        end
      end
      if((alu_write_rd_vld && (alu_write_rd_index == 5'h0d))) begin
        x_13 <= alu_write_rd_data; // @[registers.scala 79:14]
      end else begin
        if((lsu_write_normal_regfile_vld && (lsu_write_normal_rd_index == 5'h0d))) begin
          x_13 <= lsu_write_normal_rd_data; // @[registers.scala 81:14]
        end else begin
          if(lsu_write_vector_regfile_vld) begin
            if((write_vector_rd_index_0 == 5'h0d)) begin
              x_13 <= write_vector_rd_data_0; // @[registers.scala 85:18]
            end
            if((write_vector_rd_index_1 == 5'h0d)) begin
              x_13 <= write_vector_rd_data_1; // @[registers.scala 85:18]
            end
            if((write_vector_rd_index_2 == 5'h0d)) begin
              x_13 <= write_vector_rd_data_2; // @[registers.scala 85:18]
            end
            if((write_vector_rd_index_3 == 5'h0d)) begin
              x_13 <= write_vector_rd_data_3; // @[registers.scala 85:18]
            end
          end
        end
      end
      if((alu_write_rd_vld && (alu_write_rd_index == 5'h0e))) begin
        x_14 <= alu_write_rd_data; // @[registers.scala 79:14]
      end else begin
        if((lsu_write_normal_regfile_vld && (lsu_write_normal_rd_index == 5'h0e))) begin
          x_14 <= lsu_write_normal_rd_data; // @[registers.scala 81:14]
        end else begin
          if(lsu_write_vector_regfile_vld) begin
            if((write_vector_rd_index_0 == 5'h0e)) begin
              x_14 <= write_vector_rd_data_0; // @[registers.scala 85:18]
            end
            if((write_vector_rd_index_1 == 5'h0e)) begin
              x_14 <= write_vector_rd_data_1; // @[registers.scala 85:18]
            end
            if((write_vector_rd_index_2 == 5'h0e)) begin
              x_14 <= write_vector_rd_data_2; // @[registers.scala 85:18]
            end
            if((write_vector_rd_index_3 == 5'h0e)) begin
              x_14 <= write_vector_rd_data_3; // @[registers.scala 85:18]
            end
          end
        end
      end
      if((alu_write_rd_vld && (alu_write_rd_index == 5'h0f))) begin
        x_15 <= alu_write_rd_data; // @[registers.scala 79:14]
      end else begin
        if((lsu_write_normal_regfile_vld && (lsu_write_normal_rd_index == 5'h0f))) begin
          x_15 <= lsu_write_normal_rd_data; // @[registers.scala 81:14]
        end else begin
          if(lsu_write_vector_regfile_vld) begin
            if((write_vector_rd_index_0 == 5'h0f)) begin
              x_15 <= write_vector_rd_data_0; // @[registers.scala 85:18]
            end
            if((write_vector_rd_index_1 == 5'h0f)) begin
              x_15 <= write_vector_rd_data_1; // @[registers.scala 85:18]
            end
            if((write_vector_rd_index_2 == 5'h0f)) begin
              x_15 <= write_vector_rd_data_2; // @[registers.scala 85:18]
            end
            if((write_vector_rd_index_3 == 5'h0f)) begin
              x_15 <= write_vector_rd_data_3; // @[registers.scala 85:18]
            end
          end
        end
      end
      if((alu_write_rd_vld && (alu_write_rd_index == 5'h10))) begin
        x_16 <= alu_write_rd_data; // @[registers.scala 79:14]
      end else begin
        if((lsu_write_normal_regfile_vld && (lsu_write_normal_rd_index == 5'h10))) begin
          x_16 <= lsu_write_normal_rd_data; // @[registers.scala 81:14]
        end else begin
          if(lsu_write_vector_regfile_vld) begin
            if((write_vector_rd_index_0 == 5'h10)) begin
              x_16 <= write_vector_rd_data_0; // @[registers.scala 85:18]
            end
            if((write_vector_rd_index_1 == 5'h10)) begin
              x_16 <= write_vector_rd_data_1; // @[registers.scala 85:18]
            end
            if((write_vector_rd_index_2 == 5'h10)) begin
              x_16 <= write_vector_rd_data_2; // @[registers.scala 85:18]
            end
            if((write_vector_rd_index_3 == 5'h10)) begin
              x_16 <= write_vector_rd_data_3; // @[registers.scala 85:18]
            end
          end
        end
      end
      if((alu_write_rd_vld && (alu_write_rd_index == 5'h11))) begin
        x_17 <= alu_write_rd_data; // @[registers.scala 79:14]
      end else begin
        if((lsu_write_normal_regfile_vld && (lsu_write_normal_rd_index == 5'h11))) begin
          x_17 <= lsu_write_normal_rd_data; // @[registers.scala 81:14]
        end else begin
          if(lsu_write_vector_regfile_vld) begin
            if((write_vector_rd_index_0 == 5'h11)) begin
              x_17 <= write_vector_rd_data_0; // @[registers.scala 85:18]
            end
            if((write_vector_rd_index_1 == 5'h11)) begin
              x_17 <= write_vector_rd_data_1; // @[registers.scala 85:18]
            end
            if((write_vector_rd_index_2 == 5'h11)) begin
              x_17 <= write_vector_rd_data_2; // @[registers.scala 85:18]
            end
            if((write_vector_rd_index_3 == 5'h11)) begin
              x_17 <= write_vector_rd_data_3; // @[registers.scala 85:18]
            end
          end
        end
      end
      if((alu_write_rd_vld && (alu_write_rd_index == 5'h12))) begin
        x_18 <= alu_write_rd_data; // @[registers.scala 79:14]
      end else begin
        if((lsu_write_normal_regfile_vld && (lsu_write_normal_rd_index == 5'h12))) begin
          x_18 <= lsu_write_normal_rd_data; // @[registers.scala 81:14]
        end else begin
          if(lsu_write_vector_regfile_vld) begin
            if((write_vector_rd_index_0 == 5'h12)) begin
              x_18 <= write_vector_rd_data_0; // @[registers.scala 85:18]
            end
            if((write_vector_rd_index_1 == 5'h12)) begin
              x_18 <= write_vector_rd_data_1; // @[registers.scala 85:18]
            end
            if((write_vector_rd_index_2 == 5'h12)) begin
              x_18 <= write_vector_rd_data_2; // @[registers.scala 85:18]
            end
            if((write_vector_rd_index_3 == 5'h12)) begin
              x_18 <= write_vector_rd_data_3; // @[registers.scala 85:18]
            end
          end
        end
      end
      if((alu_write_rd_vld && (alu_write_rd_index == 5'h13))) begin
        x_19 <= alu_write_rd_data; // @[registers.scala 79:14]
      end else begin
        if((lsu_write_normal_regfile_vld && (lsu_write_normal_rd_index == 5'h13))) begin
          x_19 <= lsu_write_normal_rd_data; // @[registers.scala 81:14]
        end else begin
          if(lsu_write_vector_regfile_vld) begin
            if((write_vector_rd_index_0 == 5'h13)) begin
              x_19 <= write_vector_rd_data_0; // @[registers.scala 85:18]
            end
            if((write_vector_rd_index_1 == 5'h13)) begin
              x_19 <= write_vector_rd_data_1; // @[registers.scala 85:18]
            end
            if((write_vector_rd_index_2 == 5'h13)) begin
              x_19 <= write_vector_rd_data_2; // @[registers.scala 85:18]
            end
            if((write_vector_rd_index_3 == 5'h13)) begin
              x_19 <= write_vector_rd_data_3; // @[registers.scala 85:18]
            end
          end
        end
      end
      if((alu_write_rd_vld && (alu_write_rd_index == 5'h14))) begin
        x_20 <= alu_write_rd_data; // @[registers.scala 79:14]
      end else begin
        if((lsu_write_normal_regfile_vld && (lsu_write_normal_rd_index == 5'h14))) begin
          x_20 <= lsu_write_normal_rd_data; // @[registers.scala 81:14]
        end else begin
          if(lsu_write_vector_regfile_vld) begin
            if((write_vector_rd_index_0 == 5'h14)) begin
              x_20 <= write_vector_rd_data_0; // @[registers.scala 85:18]
            end
            if((write_vector_rd_index_1 == 5'h14)) begin
              x_20 <= write_vector_rd_data_1; // @[registers.scala 85:18]
            end
            if((write_vector_rd_index_2 == 5'h14)) begin
              x_20 <= write_vector_rd_data_2; // @[registers.scala 85:18]
            end
            if((write_vector_rd_index_3 == 5'h14)) begin
              x_20 <= write_vector_rd_data_3; // @[registers.scala 85:18]
            end
          end
        end
      end
      if((alu_write_rd_vld && (alu_write_rd_index == 5'h15))) begin
        x_21 <= alu_write_rd_data; // @[registers.scala 79:14]
      end else begin
        if((lsu_write_normal_regfile_vld && (lsu_write_normal_rd_index == 5'h15))) begin
          x_21 <= lsu_write_normal_rd_data; // @[registers.scala 81:14]
        end else begin
          if(lsu_write_vector_regfile_vld) begin
            if((write_vector_rd_index_0 == 5'h15)) begin
              x_21 <= write_vector_rd_data_0; // @[registers.scala 85:18]
            end
            if((write_vector_rd_index_1 == 5'h15)) begin
              x_21 <= write_vector_rd_data_1; // @[registers.scala 85:18]
            end
            if((write_vector_rd_index_2 == 5'h15)) begin
              x_21 <= write_vector_rd_data_2; // @[registers.scala 85:18]
            end
            if((write_vector_rd_index_3 == 5'h15)) begin
              x_21 <= write_vector_rd_data_3; // @[registers.scala 85:18]
            end
          end
        end
      end
      if((alu_write_rd_vld && (alu_write_rd_index == 5'h16))) begin
        x_22 <= alu_write_rd_data; // @[registers.scala 79:14]
      end else begin
        if((lsu_write_normal_regfile_vld && (lsu_write_normal_rd_index == 5'h16))) begin
          x_22 <= lsu_write_normal_rd_data; // @[registers.scala 81:14]
        end else begin
          if(lsu_write_vector_regfile_vld) begin
            if((write_vector_rd_index_0 == 5'h16)) begin
              x_22 <= write_vector_rd_data_0; // @[registers.scala 85:18]
            end
            if((write_vector_rd_index_1 == 5'h16)) begin
              x_22 <= write_vector_rd_data_1; // @[registers.scala 85:18]
            end
            if((write_vector_rd_index_2 == 5'h16)) begin
              x_22 <= write_vector_rd_data_2; // @[registers.scala 85:18]
            end
            if((write_vector_rd_index_3 == 5'h16)) begin
              x_22 <= write_vector_rd_data_3; // @[registers.scala 85:18]
            end
          end
        end
      end
      if((alu_write_rd_vld && (alu_write_rd_index == 5'h17))) begin
        x_23 <= alu_write_rd_data; // @[registers.scala 79:14]
      end else begin
        if((lsu_write_normal_regfile_vld && (lsu_write_normal_rd_index == 5'h17))) begin
          x_23 <= lsu_write_normal_rd_data; // @[registers.scala 81:14]
        end else begin
          if(lsu_write_vector_regfile_vld) begin
            if((write_vector_rd_index_0 == 5'h17)) begin
              x_23 <= write_vector_rd_data_0; // @[registers.scala 85:18]
            end
            if((write_vector_rd_index_1 == 5'h17)) begin
              x_23 <= write_vector_rd_data_1; // @[registers.scala 85:18]
            end
            if((write_vector_rd_index_2 == 5'h17)) begin
              x_23 <= write_vector_rd_data_2; // @[registers.scala 85:18]
            end
            if((write_vector_rd_index_3 == 5'h17)) begin
              x_23 <= write_vector_rd_data_3; // @[registers.scala 85:18]
            end
          end
        end
      end
      if((alu_write_rd_vld && (alu_write_rd_index == 5'h18))) begin
        x_24 <= alu_write_rd_data; // @[registers.scala 79:14]
      end else begin
        if((lsu_write_normal_regfile_vld && (lsu_write_normal_rd_index == 5'h18))) begin
          x_24 <= lsu_write_normal_rd_data; // @[registers.scala 81:14]
        end else begin
          if(lsu_write_vector_regfile_vld) begin
            if((write_vector_rd_index_0 == 5'h18)) begin
              x_24 <= write_vector_rd_data_0; // @[registers.scala 85:18]
            end
            if((write_vector_rd_index_1 == 5'h18)) begin
              x_24 <= write_vector_rd_data_1; // @[registers.scala 85:18]
            end
            if((write_vector_rd_index_2 == 5'h18)) begin
              x_24 <= write_vector_rd_data_2; // @[registers.scala 85:18]
            end
            if((write_vector_rd_index_3 == 5'h18)) begin
              x_24 <= write_vector_rd_data_3; // @[registers.scala 85:18]
            end
          end
        end
      end
      if((alu_write_rd_vld && (alu_write_rd_index == 5'h19))) begin
        x_25 <= alu_write_rd_data; // @[registers.scala 79:14]
      end else begin
        if((lsu_write_normal_regfile_vld && (lsu_write_normal_rd_index == 5'h19))) begin
          x_25 <= lsu_write_normal_rd_data; // @[registers.scala 81:14]
        end else begin
          if(lsu_write_vector_regfile_vld) begin
            if((write_vector_rd_index_0 == 5'h19)) begin
              x_25 <= write_vector_rd_data_0; // @[registers.scala 85:18]
            end
            if((write_vector_rd_index_1 == 5'h19)) begin
              x_25 <= write_vector_rd_data_1; // @[registers.scala 85:18]
            end
            if((write_vector_rd_index_2 == 5'h19)) begin
              x_25 <= write_vector_rd_data_2; // @[registers.scala 85:18]
            end
            if((write_vector_rd_index_3 == 5'h19)) begin
              x_25 <= write_vector_rd_data_3; // @[registers.scala 85:18]
            end
          end
        end
      end
      if((alu_write_rd_vld && (alu_write_rd_index == 5'h1a))) begin
        x_26 <= alu_write_rd_data; // @[registers.scala 79:14]
      end else begin
        if((lsu_write_normal_regfile_vld && (lsu_write_normal_rd_index == 5'h1a))) begin
          x_26 <= lsu_write_normal_rd_data; // @[registers.scala 81:14]
        end else begin
          if(lsu_write_vector_regfile_vld) begin
            if((write_vector_rd_index_0 == 5'h1a)) begin
              x_26 <= write_vector_rd_data_0; // @[registers.scala 85:18]
            end
            if((write_vector_rd_index_1 == 5'h1a)) begin
              x_26 <= write_vector_rd_data_1; // @[registers.scala 85:18]
            end
            if((write_vector_rd_index_2 == 5'h1a)) begin
              x_26 <= write_vector_rd_data_2; // @[registers.scala 85:18]
            end
            if((write_vector_rd_index_3 == 5'h1a)) begin
              x_26 <= write_vector_rd_data_3; // @[registers.scala 85:18]
            end
          end
        end
      end
      if((alu_write_rd_vld && (alu_write_rd_index == 5'h1b))) begin
        x_27 <= alu_write_rd_data; // @[registers.scala 79:14]
      end else begin
        if((lsu_write_normal_regfile_vld && (lsu_write_normal_rd_index == 5'h1b))) begin
          x_27 <= lsu_write_normal_rd_data; // @[registers.scala 81:14]
        end else begin
          if(lsu_write_vector_regfile_vld) begin
            if((write_vector_rd_index_0 == 5'h1b)) begin
              x_27 <= write_vector_rd_data_0; // @[registers.scala 85:18]
            end
            if((write_vector_rd_index_1 == 5'h1b)) begin
              x_27 <= write_vector_rd_data_1; // @[registers.scala 85:18]
            end
            if((write_vector_rd_index_2 == 5'h1b)) begin
              x_27 <= write_vector_rd_data_2; // @[registers.scala 85:18]
            end
            if((write_vector_rd_index_3 == 5'h1b)) begin
              x_27 <= write_vector_rd_data_3; // @[registers.scala 85:18]
            end
          end
        end
      end
      if((alu_write_rd_vld && (alu_write_rd_index == 5'h1c))) begin
        x_28 <= alu_write_rd_data; // @[registers.scala 79:14]
      end else begin
        if((lsu_write_normal_regfile_vld && (lsu_write_normal_rd_index == 5'h1c))) begin
          x_28 <= lsu_write_normal_rd_data; // @[registers.scala 81:14]
        end else begin
          if(lsu_write_vector_regfile_vld) begin
            if((write_vector_rd_index_0 == 5'h1c)) begin
              x_28 <= write_vector_rd_data_0; // @[registers.scala 85:18]
            end
            if((write_vector_rd_index_1 == 5'h1c)) begin
              x_28 <= write_vector_rd_data_1; // @[registers.scala 85:18]
            end
            if((write_vector_rd_index_2 == 5'h1c)) begin
              x_28 <= write_vector_rd_data_2; // @[registers.scala 85:18]
            end
            if((write_vector_rd_index_3 == 5'h1c)) begin
              x_28 <= write_vector_rd_data_3; // @[registers.scala 85:18]
            end
          end
        end
      end
      if((alu_write_rd_vld && (alu_write_rd_index == 5'h1d))) begin
        x_29 <= alu_write_rd_data; // @[registers.scala 79:14]
      end else begin
        if((lsu_write_normal_regfile_vld && (lsu_write_normal_rd_index == 5'h1d))) begin
          x_29 <= lsu_write_normal_rd_data; // @[registers.scala 81:14]
        end else begin
          if(lsu_write_vector_regfile_vld) begin
            if((write_vector_rd_index_0 == 5'h1d)) begin
              x_29 <= write_vector_rd_data_0; // @[registers.scala 85:18]
            end
            if((write_vector_rd_index_1 == 5'h1d)) begin
              x_29 <= write_vector_rd_data_1; // @[registers.scala 85:18]
            end
            if((write_vector_rd_index_2 == 5'h1d)) begin
              x_29 <= write_vector_rd_data_2; // @[registers.scala 85:18]
            end
            if((write_vector_rd_index_3 == 5'h1d)) begin
              x_29 <= write_vector_rd_data_3; // @[registers.scala 85:18]
            end
          end
        end
      end
      if((alu_write_rd_vld && (alu_write_rd_index == 5'h1e))) begin
        x_30 <= alu_write_rd_data; // @[registers.scala 79:14]
      end else begin
        if((lsu_write_normal_regfile_vld && (lsu_write_normal_rd_index == 5'h1e))) begin
          x_30 <= lsu_write_normal_rd_data; // @[registers.scala 81:14]
        end else begin
          if(lsu_write_vector_regfile_vld) begin
            if((write_vector_rd_index_0 == 5'h1e)) begin
              x_30 <= write_vector_rd_data_0; // @[registers.scala 85:18]
            end
            if((write_vector_rd_index_1 == 5'h1e)) begin
              x_30 <= write_vector_rd_data_1; // @[registers.scala 85:18]
            end
            if((write_vector_rd_index_2 == 5'h1e)) begin
              x_30 <= write_vector_rd_data_2; // @[registers.scala 85:18]
            end
            if((write_vector_rd_index_3 == 5'h1e)) begin
              x_30 <= write_vector_rd_data_3; // @[registers.scala 85:18]
            end
          end
        end
      end
      if((alu_write_rd_vld && (alu_write_rd_index == 5'h1f))) begin
        x_31 <= alu_write_rd_data; // @[registers.scala 79:14]
      end else begin
        if((lsu_write_normal_regfile_vld && (lsu_write_normal_rd_index == 5'h1f))) begin
          x_31 <= lsu_write_normal_rd_data; // @[registers.scala 81:14]
        end else begin
          if(lsu_write_vector_regfile_vld) begin
            if((write_vector_rd_index_0 == 5'h1f)) begin
              x_31 <= write_vector_rd_data_0; // @[registers.scala 85:18]
            end
            if((write_vector_rd_index_1 == 5'h1f)) begin
              x_31 <= write_vector_rd_data_1; // @[registers.scala 85:18]
            end
            if((write_vector_rd_index_2 == 5'h1f)) begin
              x_31 <= write_vector_rd_data_2; // @[registers.scala 85:18]
            end
            if((write_vector_rd_index_3 == 5'h1f)) begin
              x_31 <= write_vector_rd_data_3; // @[registers.scala 85:18]
            end
          end
        end
      end
    end
  end


endmodule
