// Generator : SpinalHDL v1.8.0    git head : 4e3563a282582b41f4eaafc503787757251d23ea
// Component : win_rom
// Git hash  : 85ee573ec2fdedb6c3867ea06589ef2968a1a761

`timescale 1ns/1ps 
module win_rom (
  input      [7:0]    win_addr,
  output     [7:0]    win
);

  reg        [7:0]    tmp_win;
  wire       [7:0]    win_data_0;
  wire       [7:0]    win_data_1;
  wire       [7:0]    win_data_2;
  wire       [7:0]    win_data_3;
  wire       [7:0]    win_data_4;
  wire       [7:0]    win_data_5;
  wire       [7:0]    win_data_6;
  wire       [7:0]    win_data_7;
  wire       [7:0]    win_data_8;
  wire       [7:0]    win_data_9;
  wire       [7:0]    win_data_10;
  wire       [7:0]    win_data_11;
  wire       [7:0]    win_data_12;
  wire       [7:0]    win_data_13;
  wire       [7:0]    win_data_14;
  wire       [7:0]    win_data_15;
  wire       [7:0]    win_data_16;
  wire       [7:0]    win_data_17;
  wire       [7:0]    win_data_18;
  wire       [7:0]    win_data_19;
  wire       [7:0]    win_data_20;
  wire       [7:0]    win_data_21;
  wire       [7:0]    win_data_22;
  wire       [7:0]    win_data_23;
  wire       [7:0]    win_data_24;
  wire       [7:0]    win_data_25;
  wire       [7:0]    win_data_26;
  wire       [7:0]    win_data_27;
  wire       [7:0]    win_data_28;
  wire       [7:0]    win_data_29;
  wire       [7:0]    win_data_30;
  wire       [7:0]    win_data_31;
  wire       [7:0]    win_data_32;
  wire       [7:0]    win_data_33;
  wire       [7:0]    win_data_34;
  wire       [7:0]    win_data_35;
  wire       [7:0]    win_data_36;
  wire       [7:0]    win_data_37;
  wire       [7:0]    win_data_38;
  wire       [7:0]    win_data_39;
  wire       [7:0]    win_data_40;
  wire       [7:0]    win_data_41;
  wire       [7:0]    win_data_42;
  wire       [7:0]    win_data_43;
  wire       [7:0]    win_data_44;
  wire       [7:0]    win_data_45;
  wire       [7:0]    win_data_46;
  wire       [7:0]    win_data_47;
  wire       [7:0]    win_data_48;
  wire       [7:0]    win_data_49;
  wire       [7:0]    win_data_50;
  wire       [7:0]    win_data_51;
  wire       [7:0]    win_data_52;
  wire       [7:0]    win_data_53;
  wire       [7:0]    win_data_54;
  wire       [7:0]    win_data_55;
  wire       [7:0]    win_data_56;
  wire       [7:0]    win_data_57;
  wire       [7:0]    win_data_58;
  wire       [7:0]    win_data_59;
  wire       [7:0]    win_data_60;
  wire       [7:0]    win_data_61;
  wire       [7:0]    win_data_62;
  wire       [7:0]    win_data_63;
  wire       [7:0]    win_data_64;
  wire       [7:0]    win_data_65;
  wire       [7:0]    win_data_66;
  wire       [7:0]    win_data_67;
  wire       [7:0]    win_data_68;
  wire       [7:0]    win_data_69;
  wire       [7:0]    win_data_70;
  wire       [7:0]    win_data_71;
  wire       [7:0]    win_data_72;
  wire       [7:0]    win_data_73;
  wire       [7:0]    win_data_74;
  wire       [7:0]    win_data_75;
  wire       [7:0]    win_data_76;
  wire       [7:0]    win_data_77;
  wire       [7:0]    win_data_78;
  wire       [7:0]    win_data_79;
  wire       [7:0]    win_data_80;
  wire       [7:0]    win_data_81;
  wire       [7:0]    win_data_82;
  wire       [7:0]    win_data_83;
  wire       [7:0]    win_data_84;
  wire       [7:0]    win_data_85;
  wire       [7:0]    win_data_86;
  wire       [7:0]    win_data_87;
  wire       [7:0]    win_data_88;
  wire       [7:0]    win_data_89;
  wire       [7:0]    win_data_90;
  wire       [7:0]    win_data_91;
  wire       [7:0]    win_data_92;
  wire       [7:0]    win_data_93;
  wire       [7:0]    win_data_94;
  wire       [7:0]    win_data_95;
  wire       [7:0]    win_data_96;
  wire       [7:0]    win_data_97;
  wire       [7:0]    win_data_98;
  wire       [7:0]    win_data_99;
  wire       [7:0]    win_data_100;
  wire       [7:0]    win_data_101;
  wire       [7:0]    win_data_102;
  wire       [7:0]    win_data_103;
  wire       [7:0]    win_data_104;
  wire       [7:0]    win_data_105;
  wire       [7:0]    win_data_106;
  wire       [7:0]    win_data_107;
  wire       [7:0]    win_data_108;
  wire       [7:0]    win_data_109;
  wire       [7:0]    win_data_110;
  wire       [7:0]    win_data_111;
  wire       [7:0]    win_data_112;
  wire       [7:0]    win_data_113;
  wire       [7:0]    win_data_114;
  wire       [7:0]    win_data_115;
  wire       [7:0]    win_data_116;
  wire       [7:0]    win_data_117;
  wire       [7:0]    win_data_118;
  wire       [7:0]    win_data_119;
  wire       [7:0]    win_data_120;
  wire       [7:0]    win_data_121;
  wire       [7:0]    win_data_122;
  wire       [7:0]    win_data_123;
  wire       [7:0]    win_data_124;
  wire       [7:0]    win_data_125;
  wire       [7:0]    win_data_126;
  wire       [7:0]    win_data_127;
  wire       [7:0]    win_data_128;
  wire       [7:0]    win_data_129;
  wire       [7:0]    win_data_130;
  wire       [7:0]    win_data_131;
  wire       [7:0]    win_data_132;
  wire       [7:0]    win_data_133;
  wire       [7:0]    win_data_134;
  wire       [7:0]    win_data_135;
  wire       [7:0]    win_data_136;
  wire       [7:0]    win_data_137;
  wire       [7:0]    win_data_138;
  wire       [7:0]    win_data_139;
  wire       [7:0]    win_data_140;
  wire       [7:0]    win_data_141;
  wire       [7:0]    win_data_142;
  wire       [7:0]    win_data_143;
  wire       [7:0]    win_data_144;
  wire       [7:0]    win_data_145;
  wire       [7:0]    win_data_146;
  wire       [7:0]    win_data_147;
  wire       [7:0]    win_data_148;
  wire       [7:0]    win_data_149;
  wire       [7:0]    win_data_150;
  wire       [7:0]    win_data_151;
  wire       [7:0]    win_data_152;
  wire       [7:0]    win_data_153;
  wire       [7:0]    win_data_154;
  wire       [7:0]    win_data_155;
  wire       [7:0]    win_data_156;
  wire       [7:0]    win_data_157;
  wire       [7:0]    win_data_158;
  wire       [7:0]    win_data_159;
  wire       [7:0]    win_data_160;
  wire       [7:0]    win_data_161;
  wire       [7:0]    win_data_162;
  wire       [7:0]    win_data_163;
  wire       [7:0]    win_data_164;
  wire       [7:0]    win_data_165;
  wire       [7:0]    win_data_166;
  wire       [7:0]    win_data_167;
  wire       [7:0]    win_data_168;
  wire       [7:0]    win_data_169;
  wire       [7:0]    win_data_170;
  wire       [7:0]    win_data_171;
  wire       [7:0]    win_data_172;
  wire       [7:0]    win_data_173;
  wire       [7:0]    win_data_174;
  wire       [7:0]    win_data_175;
  wire       [7:0]    win_data_176;
  wire       [7:0]    win_data_177;
  wire       [7:0]    win_data_178;
  wire       [7:0]    win_data_179;
  wire       [7:0]    win_data_180;
  wire       [7:0]    win_data_181;
  wire       [7:0]    win_data_182;
  wire       [7:0]    win_data_183;
  wire       [7:0]    win_data_184;
  wire       [7:0]    win_data_185;
  wire       [7:0]    win_data_186;
  wire       [7:0]    win_data_187;
  wire       [7:0]    win_data_188;
  wire       [7:0]    win_data_189;
  wire       [7:0]    win_data_190;
  wire       [7:0]    win_data_191;
  wire       [7:0]    win_data_192;
  wire       [7:0]    win_data_193;
  wire       [7:0]    win_data_194;
  wire       [7:0]    win_data_195;
  wire       [7:0]    win_data_196;
  wire       [7:0]    win_data_197;
  wire       [7:0]    win_data_198;
  wire       [7:0]    win_data_199;
  wire       [7:0]    win_data_200;
  wire       [7:0]    win_data_201;
  wire       [7:0]    win_data_202;
  wire       [7:0]    win_data_203;
  wire       [7:0]    win_data_204;
  wire       [7:0]    win_data_205;
  wire       [7:0]    win_data_206;
  wire       [7:0]    win_data_207;
  wire       [7:0]    win_data_208;
  wire       [7:0]    win_data_209;
  wire       [7:0]    win_data_210;
  wire       [7:0]    win_data_211;
  wire       [7:0]    win_data_212;
  wire       [7:0]    win_data_213;
  wire       [7:0]    win_data_214;
  wire       [7:0]    win_data_215;
  wire       [7:0]    win_data_216;
  wire       [7:0]    win_data_217;
  wire       [7:0]    win_data_218;
  wire       [7:0]    win_data_219;
  wire       [7:0]    win_data_220;
  wire       [7:0]    win_data_221;
  wire       [7:0]    win_data_222;
  wire       [7:0]    win_data_223;
  wire       [7:0]    win_data_224;
  wire       [7:0]    win_data_225;
  wire       [7:0]    win_data_226;
  wire       [7:0]    win_data_227;
  wire       [7:0]    win_data_228;
  wire       [7:0]    win_data_229;
  wire       [7:0]    win_data_230;
  wire       [7:0]    win_data_231;
  wire       [7:0]    win_data_232;
  wire       [7:0]    win_data_233;
  wire       [7:0]    win_data_234;
  wire       [7:0]    win_data_235;
  wire       [7:0]    win_data_236;
  wire       [7:0]    win_data_237;
  wire       [7:0]    win_data_238;
  wire       [7:0]    win_data_239;
  wire       [7:0]    win_data_240;
  wire       [7:0]    win_data_241;
  wire       [7:0]    win_data_242;
  wire       [7:0]    win_data_243;
  wire       [7:0]    win_data_244;
  wire       [7:0]    win_data_245;
  wire       [7:0]    win_data_246;
  wire       [7:0]    win_data_247;
  wire       [7:0]    win_data_248;
  wire       [7:0]    win_data_249;
  wire       [7:0]    win_data_250;
  wire       [7:0]    win_data_251;
  wire       [7:0]    win_data_252;
  wire       [7:0]    win_data_253;
  wire       [7:0]    win_data_254;
  wire       [7:0]    win_data_255;

  always @(*) begin
    case(win_addr)
      8'b00000000 : tmp_win = win_data_0;
      8'b00000001 : tmp_win = win_data_1;
      8'b00000010 : tmp_win = win_data_2;
      8'b00000011 : tmp_win = win_data_3;
      8'b00000100 : tmp_win = win_data_4;
      8'b00000101 : tmp_win = win_data_5;
      8'b00000110 : tmp_win = win_data_6;
      8'b00000111 : tmp_win = win_data_7;
      8'b00001000 : tmp_win = win_data_8;
      8'b00001001 : tmp_win = win_data_9;
      8'b00001010 : tmp_win = win_data_10;
      8'b00001011 : tmp_win = win_data_11;
      8'b00001100 : tmp_win = win_data_12;
      8'b00001101 : tmp_win = win_data_13;
      8'b00001110 : tmp_win = win_data_14;
      8'b00001111 : tmp_win = win_data_15;
      8'b00010000 : tmp_win = win_data_16;
      8'b00010001 : tmp_win = win_data_17;
      8'b00010010 : tmp_win = win_data_18;
      8'b00010011 : tmp_win = win_data_19;
      8'b00010100 : tmp_win = win_data_20;
      8'b00010101 : tmp_win = win_data_21;
      8'b00010110 : tmp_win = win_data_22;
      8'b00010111 : tmp_win = win_data_23;
      8'b00011000 : tmp_win = win_data_24;
      8'b00011001 : tmp_win = win_data_25;
      8'b00011010 : tmp_win = win_data_26;
      8'b00011011 : tmp_win = win_data_27;
      8'b00011100 : tmp_win = win_data_28;
      8'b00011101 : tmp_win = win_data_29;
      8'b00011110 : tmp_win = win_data_30;
      8'b00011111 : tmp_win = win_data_31;
      8'b00100000 : tmp_win = win_data_32;
      8'b00100001 : tmp_win = win_data_33;
      8'b00100010 : tmp_win = win_data_34;
      8'b00100011 : tmp_win = win_data_35;
      8'b00100100 : tmp_win = win_data_36;
      8'b00100101 : tmp_win = win_data_37;
      8'b00100110 : tmp_win = win_data_38;
      8'b00100111 : tmp_win = win_data_39;
      8'b00101000 : tmp_win = win_data_40;
      8'b00101001 : tmp_win = win_data_41;
      8'b00101010 : tmp_win = win_data_42;
      8'b00101011 : tmp_win = win_data_43;
      8'b00101100 : tmp_win = win_data_44;
      8'b00101101 : tmp_win = win_data_45;
      8'b00101110 : tmp_win = win_data_46;
      8'b00101111 : tmp_win = win_data_47;
      8'b00110000 : tmp_win = win_data_48;
      8'b00110001 : tmp_win = win_data_49;
      8'b00110010 : tmp_win = win_data_50;
      8'b00110011 : tmp_win = win_data_51;
      8'b00110100 : tmp_win = win_data_52;
      8'b00110101 : tmp_win = win_data_53;
      8'b00110110 : tmp_win = win_data_54;
      8'b00110111 : tmp_win = win_data_55;
      8'b00111000 : tmp_win = win_data_56;
      8'b00111001 : tmp_win = win_data_57;
      8'b00111010 : tmp_win = win_data_58;
      8'b00111011 : tmp_win = win_data_59;
      8'b00111100 : tmp_win = win_data_60;
      8'b00111101 : tmp_win = win_data_61;
      8'b00111110 : tmp_win = win_data_62;
      8'b00111111 : tmp_win = win_data_63;
      8'b01000000 : tmp_win = win_data_64;
      8'b01000001 : tmp_win = win_data_65;
      8'b01000010 : tmp_win = win_data_66;
      8'b01000011 : tmp_win = win_data_67;
      8'b01000100 : tmp_win = win_data_68;
      8'b01000101 : tmp_win = win_data_69;
      8'b01000110 : tmp_win = win_data_70;
      8'b01000111 : tmp_win = win_data_71;
      8'b01001000 : tmp_win = win_data_72;
      8'b01001001 : tmp_win = win_data_73;
      8'b01001010 : tmp_win = win_data_74;
      8'b01001011 : tmp_win = win_data_75;
      8'b01001100 : tmp_win = win_data_76;
      8'b01001101 : tmp_win = win_data_77;
      8'b01001110 : tmp_win = win_data_78;
      8'b01001111 : tmp_win = win_data_79;
      8'b01010000 : tmp_win = win_data_80;
      8'b01010001 : tmp_win = win_data_81;
      8'b01010010 : tmp_win = win_data_82;
      8'b01010011 : tmp_win = win_data_83;
      8'b01010100 : tmp_win = win_data_84;
      8'b01010101 : tmp_win = win_data_85;
      8'b01010110 : tmp_win = win_data_86;
      8'b01010111 : tmp_win = win_data_87;
      8'b01011000 : tmp_win = win_data_88;
      8'b01011001 : tmp_win = win_data_89;
      8'b01011010 : tmp_win = win_data_90;
      8'b01011011 : tmp_win = win_data_91;
      8'b01011100 : tmp_win = win_data_92;
      8'b01011101 : tmp_win = win_data_93;
      8'b01011110 : tmp_win = win_data_94;
      8'b01011111 : tmp_win = win_data_95;
      8'b01100000 : tmp_win = win_data_96;
      8'b01100001 : tmp_win = win_data_97;
      8'b01100010 : tmp_win = win_data_98;
      8'b01100011 : tmp_win = win_data_99;
      8'b01100100 : tmp_win = win_data_100;
      8'b01100101 : tmp_win = win_data_101;
      8'b01100110 : tmp_win = win_data_102;
      8'b01100111 : tmp_win = win_data_103;
      8'b01101000 : tmp_win = win_data_104;
      8'b01101001 : tmp_win = win_data_105;
      8'b01101010 : tmp_win = win_data_106;
      8'b01101011 : tmp_win = win_data_107;
      8'b01101100 : tmp_win = win_data_108;
      8'b01101101 : tmp_win = win_data_109;
      8'b01101110 : tmp_win = win_data_110;
      8'b01101111 : tmp_win = win_data_111;
      8'b01110000 : tmp_win = win_data_112;
      8'b01110001 : tmp_win = win_data_113;
      8'b01110010 : tmp_win = win_data_114;
      8'b01110011 : tmp_win = win_data_115;
      8'b01110100 : tmp_win = win_data_116;
      8'b01110101 : tmp_win = win_data_117;
      8'b01110110 : tmp_win = win_data_118;
      8'b01110111 : tmp_win = win_data_119;
      8'b01111000 : tmp_win = win_data_120;
      8'b01111001 : tmp_win = win_data_121;
      8'b01111010 : tmp_win = win_data_122;
      8'b01111011 : tmp_win = win_data_123;
      8'b01111100 : tmp_win = win_data_124;
      8'b01111101 : tmp_win = win_data_125;
      8'b01111110 : tmp_win = win_data_126;
      8'b01111111 : tmp_win = win_data_127;
      8'b10000000 : tmp_win = win_data_128;
      8'b10000001 : tmp_win = win_data_129;
      8'b10000010 : tmp_win = win_data_130;
      8'b10000011 : tmp_win = win_data_131;
      8'b10000100 : tmp_win = win_data_132;
      8'b10000101 : tmp_win = win_data_133;
      8'b10000110 : tmp_win = win_data_134;
      8'b10000111 : tmp_win = win_data_135;
      8'b10001000 : tmp_win = win_data_136;
      8'b10001001 : tmp_win = win_data_137;
      8'b10001010 : tmp_win = win_data_138;
      8'b10001011 : tmp_win = win_data_139;
      8'b10001100 : tmp_win = win_data_140;
      8'b10001101 : tmp_win = win_data_141;
      8'b10001110 : tmp_win = win_data_142;
      8'b10001111 : tmp_win = win_data_143;
      8'b10010000 : tmp_win = win_data_144;
      8'b10010001 : tmp_win = win_data_145;
      8'b10010010 : tmp_win = win_data_146;
      8'b10010011 : tmp_win = win_data_147;
      8'b10010100 : tmp_win = win_data_148;
      8'b10010101 : tmp_win = win_data_149;
      8'b10010110 : tmp_win = win_data_150;
      8'b10010111 : tmp_win = win_data_151;
      8'b10011000 : tmp_win = win_data_152;
      8'b10011001 : tmp_win = win_data_153;
      8'b10011010 : tmp_win = win_data_154;
      8'b10011011 : tmp_win = win_data_155;
      8'b10011100 : tmp_win = win_data_156;
      8'b10011101 : tmp_win = win_data_157;
      8'b10011110 : tmp_win = win_data_158;
      8'b10011111 : tmp_win = win_data_159;
      8'b10100000 : tmp_win = win_data_160;
      8'b10100001 : tmp_win = win_data_161;
      8'b10100010 : tmp_win = win_data_162;
      8'b10100011 : tmp_win = win_data_163;
      8'b10100100 : tmp_win = win_data_164;
      8'b10100101 : tmp_win = win_data_165;
      8'b10100110 : tmp_win = win_data_166;
      8'b10100111 : tmp_win = win_data_167;
      8'b10101000 : tmp_win = win_data_168;
      8'b10101001 : tmp_win = win_data_169;
      8'b10101010 : tmp_win = win_data_170;
      8'b10101011 : tmp_win = win_data_171;
      8'b10101100 : tmp_win = win_data_172;
      8'b10101101 : tmp_win = win_data_173;
      8'b10101110 : tmp_win = win_data_174;
      8'b10101111 : tmp_win = win_data_175;
      8'b10110000 : tmp_win = win_data_176;
      8'b10110001 : tmp_win = win_data_177;
      8'b10110010 : tmp_win = win_data_178;
      8'b10110011 : tmp_win = win_data_179;
      8'b10110100 : tmp_win = win_data_180;
      8'b10110101 : tmp_win = win_data_181;
      8'b10110110 : tmp_win = win_data_182;
      8'b10110111 : tmp_win = win_data_183;
      8'b10111000 : tmp_win = win_data_184;
      8'b10111001 : tmp_win = win_data_185;
      8'b10111010 : tmp_win = win_data_186;
      8'b10111011 : tmp_win = win_data_187;
      8'b10111100 : tmp_win = win_data_188;
      8'b10111101 : tmp_win = win_data_189;
      8'b10111110 : tmp_win = win_data_190;
      8'b10111111 : tmp_win = win_data_191;
      8'b11000000 : tmp_win = win_data_192;
      8'b11000001 : tmp_win = win_data_193;
      8'b11000010 : tmp_win = win_data_194;
      8'b11000011 : tmp_win = win_data_195;
      8'b11000100 : tmp_win = win_data_196;
      8'b11000101 : tmp_win = win_data_197;
      8'b11000110 : tmp_win = win_data_198;
      8'b11000111 : tmp_win = win_data_199;
      8'b11001000 : tmp_win = win_data_200;
      8'b11001001 : tmp_win = win_data_201;
      8'b11001010 : tmp_win = win_data_202;
      8'b11001011 : tmp_win = win_data_203;
      8'b11001100 : tmp_win = win_data_204;
      8'b11001101 : tmp_win = win_data_205;
      8'b11001110 : tmp_win = win_data_206;
      8'b11001111 : tmp_win = win_data_207;
      8'b11010000 : tmp_win = win_data_208;
      8'b11010001 : tmp_win = win_data_209;
      8'b11010010 : tmp_win = win_data_210;
      8'b11010011 : tmp_win = win_data_211;
      8'b11010100 : tmp_win = win_data_212;
      8'b11010101 : tmp_win = win_data_213;
      8'b11010110 : tmp_win = win_data_214;
      8'b11010111 : tmp_win = win_data_215;
      8'b11011000 : tmp_win = win_data_216;
      8'b11011001 : tmp_win = win_data_217;
      8'b11011010 : tmp_win = win_data_218;
      8'b11011011 : tmp_win = win_data_219;
      8'b11011100 : tmp_win = win_data_220;
      8'b11011101 : tmp_win = win_data_221;
      8'b11011110 : tmp_win = win_data_222;
      8'b11011111 : tmp_win = win_data_223;
      8'b11100000 : tmp_win = win_data_224;
      8'b11100001 : tmp_win = win_data_225;
      8'b11100010 : tmp_win = win_data_226;
      8'b11100011 : tmp_win = win_data_227;
      8'b11100100 : tmp_win = win_data_228;
      8'b11100101 : tmp_win = win_data_229;
      8'b11100110 : tmp_win = win_data_230;
      8'b11100111 : tmp_win = win_data_231;
      8'b11101000 : tmp_win = win_data_232;
      8'b11101001 : tmp_win = win_data_233;
      8'b11101010 : tmp_win = win_data_234;
      8'b11101011 : tmp_win = win_data_235;
      8'b11101100 : tmp_win = win_data_236;
      8'b11101101 : tmp_win = win_data_237;
      8'b11101110 : tmp_win = win_data_238;
      8'b11101111 : tmp_win = win_data_239;
      8'b11110000 : tmp_win = win_data_240;
      8'b11110001 : tmp_win = win_data_241;
      8'b11110010 : tmp_win = win_data_242;
      8'b11110011 : tmp_win = win_data_243;
      8'b11110100 : tmp_win = win_data_244;
      8'b11110101 : tmp_win = win_data_245;
      8'b11110110 : tmp_win = win_data_246;
      8'b11110111 : tmp_win = win_data_247;
      8'b11111000 : tmp_win = win_data_248;
      8'b11111001 : tmp_win = win_data_249;
      8'b11111010 : tmp_win = win_data_250;
      8'b11111011 : tmp_win = win_data_251;
      8'b11111100 : tmp_win = win_data_252;
      8'b11111101 : tmp_win = win_data_253;
      8'b11111110 : tmp_win = win_data_254;
      default : tmp_win = win_data_255;
    endcase
  end

  assign win_data_0 = 8'h0; // @[Expression.scala 2342:18]
  assign win_data_1 = 8'h0; // @[Expression.scala 2342:18]
  assign win_data_2 = 8'h0; // @[Expression.scala 2342:18]
  assign win_data_3 = 8'h0; // @[Expression.scala 2342:18]
  assign win_data_4 = 8'h01; // @[Expression.scala 2342:18]
  assign win_data_5 = 8'h01; // @[Expression.scala 2342:18]
  assign win_data_6 = 8'h01; // @[Expression.scala 2342:18]
  assign win_data_7 = 8'h02; // @[Expression.scala 2342:18]
  assign win_data_8 = 8'h02; // @[Expression.scala 2342:18]
  assign win_data_9 = 8'h03; // @[Expression.scala 2342:18]
  assign win_data_10 = 8'h04; // @[Expression.scala 2342:18]
  assign win_data_11 = 8'h05; // @[Expression.scala 2342:18]
  assign win_data_12 = 8'h05; // @[Expression.scala 2342:18]
  assign win_data_13 = 8'h06; // @[Expression.scala 2342:18]
  assign win_data_14 = 8'h07; // @[Expression.scala 2342:18]
  assign win_data_15 = 8'h09; // @[Expression.scala 2342:18]
  assign win_data_16 = 8'h0a; // @[Expression.scala 2342:18]
  assign win_data_17 = 8'h0b; // @[Expression.scala 2342:18]
  assign win_data_18 = 8'h0c; // @[Expression.scala 2342:18]
  assign win_data_19 = 8'h0e; // @[Expression.scala 2342:18]
  assign win_data_20 = 8'h0f; // @[Expression.scala 2342:18]
  assign win_data_21 = 8'h11; // @[Expression.scala 2342:18]
  assign win_data_22 = 8'h12; // @[Expression.scala 2342:18]
  assign win_data_23 = 8'h14; // @[Expression.scala 2342:18]
  assign win_data_24 = 8'h15; // @[Expression.scala 2342:18]
  assign win_data_25 = 8'h17; // @[Expression.scala 2342:18]
  assign win_data_26 = 8'h19; // @[Expression.scala 2342:18]
  assign win_data_27 = 8'h1b; // @[Expression.scala 2342:18]
  assign win_data_28 = 8'h1d; // @[Expression.scala 2342:18]
  assign win_data_29 = 8'h1f; // @[Expression.scala 2342:18]
  assign win_data_30 = 8'h21; // @[Expression.scala 2342:18]
  assign win_data_31 = 8'h23; // @[Expression.scala 2342:18]
  assign win_data_32 = 8'h25; // @[Expression.scala 2342:18]
  assign win_data_33 = 8'h28; // @[Expression.scala 2342:18]
  assign win_data_34 = 8'h2a; // @[Expression.scala 2342:18]
  assign win_data_35 = 8'h2c; // @[Expression.scala 2342:18]
  assign win_data_36 = 8'h2f; // @[Expression.scala 2342:18]
  assign win_data_37 = 8'h31; // @[Expression.scala 2342:18]
  assign win_data_38 = 8'h34; // @[Expression.scala 2342:18]
  assign win_data_39 = 8'h36; // @[Expression.scala 2342:18]
  assign win_data_40 = 8'h39; // @[Expression.scala 2342:18]
  assign win_data_41 = 8'h3b; // @[Expression.scala 2342:18]
  assign win_data_42 = 8'h3e; // @[Expression.scala 2342:18]
  assign win_data_43 = 8'h41; // @[Expression.scala 2342:18]
  assign win_data_44 = 8'h43; // @[Expression.scala 2342:18]
  assign win_data_45 = 8'h46; // @[Expression.scala 2342:18]
  assign win_data_46 = 8'h49; // @[Expression.scala 2342:18]
  assign win_data_47 = 8'h4c; // @[Expression.scala 2342:18]
  assign win_data_48 = 8'h4f; // @[Expression.scala 2342:18]
  assign win_data_49 = 8'h52; // @[Expression.scala 2342:18]
  assign win_data_50 = 8'h55; // @[Expression.scala 2342:18]
  assign win_data_51 = 8'h58; // @[Expression.scala 2342:18]
  assign win_data_52 = 8'h5a; // @[Expression.scala 2342:18]
  assign win_data_53 = 8'h5d; // @[Expression.scala 2342:18]
  assign win_data_54 = 8'h61; // @[Expression.scala 2342:18]
  assign win_data_55 = 8'h64; // @[Expression.scala 2342:18]
  assign win_data_56 = 8'h67; // @[Expression.scala 2342:18]
  assign win_data_57 = 8'h6a; // @[Expression.scala 2342:18]
  assign win_data_58 = 8'h6d; // @[Expression.scala 2342:18]
  assign win_data_59 = 8'h70; // @[Expression.scala 2342:18]
  assign win_data_60 = 8'h73; // @[Expression.scala 2342:18]
  assign win_data_61 = 8'h76; // @[Expression.scala 2342:18]
  assign win_data_62 = 8'h79; // @[Expression.scala 2342:18]
  assign win_data_63 = 8'h7c; // @[Expression.scala 2342:18]
  assign win_data_64 = 8'h80; // @[Expression.scala 2342:18]
  assign win_data_65 = 8'h83; // @[Expression.scala 2342:18]
  assign win_data_66 = 8'h86; // @[Expression.scala 2342:18]
  assign win_data_67 = 8'h89; // @[Expression.scala 2342:18]
  assign win_data_68 = 8'h8c; // @[Expression.scala 2342:18]
  assign win_data_69 = 8'h8f; // @[Expression.scala 2342:18]
  assign win_data_70 = 8'h92; // @[Expression.scala 2342:18]
  assign win_data_71 = 8'h95; // @[Expression.scala 2342:18]
  assign win_data_72 = 8'h98; // @[Expression.scala 2342:18]
  assign win_data_73 = 8'h9b; // @[Expression.scala 2342:18]
  assign win_data_74 = 8'h9e; // @[Expression.scala 2342:18]
  assign win_data_75 = 8'ha2; // @[Expression.scala 2342:18]
  assign win_data_76 = 8'ha5; // @[Expression.scala 2342:18]
  assign win_data_77 = 8'ha7; // @[Expression.scala 2342:18]
  assign win_data_78 = 8'haa; // @[Expression.scala 2342:18]
  assign win_data_79 = 8'had; // @[Expression.scala 2342:18]
  assign win_data_80 = 8'hb0; // @[Expression.scala 2342:18]
  assign win_data_81 = 8'hb3; // @[Expression.scala 2342:18]
  assign win_data_82 = 8'hb6; // @[Expression.scala 2342:18]
  assign win_data_83 = 8'hb9; // @[Expression.scala 2342:18]
  assign win_data_84 = 8'hbc; // @[Expression.scala 2342:18]
  assign win_data_85 = 8'hbe; // @[Expression.scala 2342:18]
  assign win_data_86 = 8'hc1; // @[Expression.scala 2342:18]
  assign win_data_87 = 8'hc4; // @[Expression.scala 2342:18]
  assign win_data_88 = 8'hc6; // @[Expression.scala 2342:18]
  assign win_data_89 = 8'hc9; // @[Expression.scala 2342:18]
  assign win_data_90 = 8'hcb; // @[Expression.scala 2342:18]
  assign win_data_91 = 8'hce; // @[Expression.scala 2342:18]
  assign win_data_92 = 8'hd0; // @[Expression.scala 2342:18]
  assign win_data_93 = 8'hd3; // @[Expression.scala 2342:18]
  assign win_data_94 = 8'hd5; // @[Expression.scala 2342:18]
  assign win_data_95 = 8'hd7; // @[Expression.scala 2342:18]
  assign win_data_96 = 8'hda; // @[Expression.scala 2342:18]
  assign win_data_97 = 8'hdc; // @[Expression.scala 2342:18]
  assign win_data_98 = 8'hde; // @[Expression.scala 2342:18]
  assign win_data_99 = 8'he0; // @[Expression.scala 2342:18]
  assign win_data_100 = 8'he2; // @[Expression.scala 2342:18]
  assign win_data_101 = 8'he4; // @[Expression.scala 2342:18]
  assign win_data_102 = 8'he6; // @[Expression.scala 2342:18]
  assign win_data_103 = 8'he8; // @[Expression.scala 2342:18]
  assign win_data_104 = 8'hea; // @[Expression.scala 2342:18]
  assign win_data_105 = 8'heb; // @[Expression.scala 2342:18]
  assign win_data_106 = 8'hed; // @[Expression.scala 2342:18]
  assign win_data_107 = 8'hee; // @[Expression.scala 2342:18]
  assign win_data_108 = 8'hf0; // @[Expression.scala 2342:18]
  assign win_data_109 = 8'hf1; // @[Expression.scala 2342:18]
  assign win_data_110 = 8'hf3; // @[Expression.scala 2342:18]
  assign win_data_111 = 8'hf4; // @[Expression.scala 2342:18]
  assign win_data_112 = 8'hf5; // @[Expression.scala 2342:18]
  assign win_data_113 = 8'hf6; // @[Expression.scala 2342:18]
  assign win_data_114 = 8'hf8; // @[Expression.scala 2342:18]
  assign win_data_115 = 8'hf9; // @[Expression.scala 2342:18]
  assign win_data_116 = 8'hfa; // @[Expression.scala 2342:18]
  assign win_data_117 = 8'hfa; // @[Expression.scala 2342:18]
  assign win_data_118 = 8'hfb; // @[Expression.scala 2342:18]
  assign win_data_119 = 8'hfc; // @[Expression.scala 2342:18]
  assign win_data_120 = 8'hfd; // @[Expression.scala 2342:18]
  assign win_data_121 = 8'hfd; // @[Expression.scala 2342:18]
  assign win_data_122 = 8'hfe; // @[Expression.scala 2342:18]
  assign win_data_123 = 8'hfe; // @[Expression.scala 2342:18]
  assign win_data_124 = 8'hfe; // @[Expression.scala 2342:18]
  assign win_data_125 = 8'hff; // @[Expression.scala 2342:18]
  assign win_data_126 = 8'hff; // @[Expression.scala 2342:18]
  assign win_data_127 = 8'hff; // @[Expression.scala 2342:18]
  assign win_data_128 = 8'hff; // @[Expression.scala 2342:18]
  assign win_data_129 = 8'hff; // @[Expression.scala 2342:18]
  assign win_data_130 = 8'hff; // @[Expression.scala 2342:18]
  assign win_data_131 = 8'hff; // @[Expression.scala 2342:18]
  assign win_data_132 = 8'hfe; // @[Expression.scala 2342:18]
  assign win_data_133 = 8'hfe; // @[Expression.scala 2342:18]
  assign win_data_134 = 8'hfe; // @[Expression.scala 2342:18]
  assign win_data_135 = 8'hfd; // @[Expression.scala 2342:18]
  assign win_data_136 = 8'hfd; // @[Expression.scala 2342:18]
  assign win_data_137 = 8'hfc; // @[Expression.scala 2342:18]
  assign win_data_138 = 8'hfb; // @[Expression.scala 2342:18]
  assign win_data_139 = 8'hfa; // @[Expression.scala 2342:18]
  assign win_data_140 = 8'hfa; // @[Expression.scala 2342:18]
  assign win_data_141 = 8'hf9; // @[Expression.scala 2342:18]
  assign win_data_142 = 8'hf8; // @[Expression.scala 2342:18]
  assign win_data_143 = 8'hf6; // @[Expression.scala 2342:18]
  assign win_data_144 = 8'hf5; // @[Expression.scala 2342:18]
  assign win_data_145 = 8'hf4; // @[Expression.scala 2342:18]
  assign win_data_146 = 8'hf3; // @[Expression.scala 2342:18]
  assign win_data_147 = 8'hf1; // @[Expression.scala 2342:18]
  assign win_data_148 = 8'hf0; // @[Expression.scala 2342:18]
  assign win_data_149 = 8'hee; // @[Expression.scala 2342:18]
  assign win_data_150 = 8'hed; // @[Expression.scala 2342:18]
  assign win_data_151 = 8'heb; // @[Expression.scala 2342:18]
  assign win_data_152 = 8'hea; // @[Expression.scala 2342:18]
  assign win_data_153 = 8'he8; // @[Expression.scala 2342:18]
  assign win_data_154 = 8'he6; // @[Expression.scala 2342:18]
  assign win_data_155 = 8'he4; // @[Expression.scala 2342:18]
  assign win_data_156 = 8'he2; // @[Expression.scala 2342:18]
  assign win_data_157 = 8'he0; // @[Expression.scala 2342:18]
  assign win_data_158 = 8'hde; // @[Expression.scala 2342:18]
  assign win_data_159 = 8'hdc; // @[Expression.scala 2342:18]
  assign win_data_160 = 8'hda; // @[Expression.scala 2342:18]
  assign win_data_161 = 8'hd7; // @[Expression.scala 2342:18]
  assign win_data_162 = 8'hd5; // @[Expression.scala 2342:18]
  assign win_data_163 = 8'hd3; // @[Expression.scala 2342:18]
  assign win_data_164 = 8'hd0; // @[Expression.scala 2342:18]
  assign win_data_165 = 8'hce; // @[Expression.scala 2342:18]
  assign win_data_166 = 8'hcb; // @[Expression.scala 2342:18]
  assign win_data_167 = 8'hc9; // @[Expression.scala 2342:18]
  assign win_data_168 = 8'hc6; // @[Expression.scala 2342:18]
  assign win_data_169 = 8'hc4; // @[Expression.scala 2342:18]
  assign win_data_170 = 8'hc1; // @[Expression.scala 2342:18]
  assign win_data_171 = 8'hbe; // @[Expression.scala 2342:18]
  assign win_data_172 = 8'hbc; // @[Expression.scala 2342:18]
  assign win_data_173 = 8'hb9; // @[Expression.scala 2342:18]
  assign win_data_174 = 8'hb6; // @[Expression.scala 2342:18]
  assign win_data_175 = 8'hb3; // @[Expression.scala 2342:18]
  assign win_data_176 = 8'hb0; // @[Expression.scala 2342:18]
  assign win_data_177 = 8'had; // @[Expression.scala 2342:18]
  assign win_data_178 = 8'haa; // @[Expression.scala 2342:18]
  assign win_data_179 = 8'ha7; // @[Expression.scala 2342:18]
  assign win_data_180 = 8'ha5; // @[Expression.scala 2342:18]
  assign win_data_181 = 8'ha2; // @[Expression.scala 2342:18]
  assign win_data_182 = 8'h9e; // @[Expression.scala 2342:18]
  assign win_data_183 = 8'h9b; // @[Expression.scala 2342:18]
  assign win_data_184 = 8'h98; // @[Expression.scala 2342:18]
  assign win_data_185 = 8'h95; // @[Expression.scala 2342:18]
  assign win_data_186 = 8'h92; // @[Expression.scala 2342:18]
  assign win_data_187 = 8'h8f; // @[Expression.scala 2342:18]
  assign win_data_188 = 8'h8c; // @[Expression.scala 2342:18]
  assign win_data_189 = 8'h89; // @[Expression.scala 2342:18]
  assign win_data_190 = 8'h86; // @[Expression.scala 2342:18]
  assign win_data_191 = 8'h83; // @[Expression.scala 2342:18]
  assign win_data_192 = 8'h80; // @[Expression.scala 2342:18]
  assign win_data_193 = 8'h7c; // @[Expression.scala 2342:18]
  assign win_data_194 = 8'h79; // @[Expression.scala 2342:18]
  assign win_data_195 = 8'h76; // @[Expression.scala 2342:18]
  assign win_data_196 = 8'h73; // @[Expression.scala 2342:18]
  assign win_data_197 = 8'h70; // @[Expression.scala 2342:18]
  assign win_data_198 = 8'h6d; // @[Expression.scala 2342:18]
  assign win_data_199 = 8'h6a; // @[Expression.scala 2342:18]
  assign win_data_200 = 8'h67; // @[Expression.scala 2342:18]
  assign win_data_201 = 8'h64; // @[Expression.scala 2342:18]
  assign win_data_202 = 8'h61; // @[Expression.scala 2342:18]
  assign win_data_203 = 8'h5d; // @[Expression.scala 2342:18]
  assign win_data_204 = 8'h5a; // @[Expression.scala 2342:18]
  assign win_data_205 = 8'h58; // @[Expression.scala 2342:18]
  assign win_data_206 = 8'h55; // @[Expression.scala 2342:18]
  assign win_data_207 = 8'h52; // @[Expression.scala 2342:18]
  assign win_data_208 = 8'h4f; // @[Expression.scala 2342:18]
  assign win_data_209 = 8'h4c; // @[Expression.scala 2342:18]
  assign win_data_210 = 8'h49; // @[Expression.scala 2342:18]
  assign win_data_211 = 8'h46; // @[Expression.scala 2342:18]
  assign win_data_212 = 8'h43; // @[Expression.scala 2342:18]
  assign win_data_213 = 8'h41; // @[Expression.scala 2342:18]
  assign win_data_214 = 8'h3e; // @[Expression.scala 2342:18]
  assign win_data_215 = 8'h3b; // @[Expression.scala 2342:18]
  assign win_data_216 = 8'h39; // @[Expression.scala 2342:18]
  assign win_data_217 = 8'h36; // @[Expression.scala 2342:18]
  assign win_data_218 = 8'h34; // @[Expression.scala 2342:18]
  assign win_data_219 = 8'h31; // @[Expression.scala 2342:18]
  assign win_data_220 = 8'h2f; // @[Expression.scala 2342:18]
  assign win_data_221 = 8'h2c; // @[Expression.scala 2342:18]
  assign win_data_222 = 8'h2a; // @[Expression.scala 2342:18]
  assign win_data_223 = 8'h28; // @[Expression.scala 2342:18]
  assign win_data_224 = 8'h25; // @[Expression.scala 2342:18]
  assign win_data_225 = 8'h23; // @[Expression.scala 2342:18]
  assign win_data_226 = 8'h21; // @[Expression.scala 2342:18]
  assign win_data_227 = 8'h1f; // @[Expression.scala 2342:18]
  assign win_data_228 = 8'h1d; // @[Expression.scala 2342:18]
  assign win_data_229 = 8'h1b; // @[Expression.scala 2342:18]
  assign win_data_230 = 8'h19; // @[Expression.scala 2342:18]
  assign win_data_231 = 8'h17; // @[Expression.scala 2342:18]
  assign win_data_232 = 8'h15; // @[Expression.scala 2342:18]
  assign win_data_233 = 8'h14; // @[Expression.scala 2342:18]
  assign win_data_234 = 8'h12; // @[Expression.scala 2342:18]
  assign win_data_235 = 8'h11; // @[Expression.scala 2342:18]
  assign win_data_236 = 8'h0f; // @[Expression.scala 2342:18]
  assign win_data_237 = 8'h0e; // @[Expression.scala 2342:18]
  assign win_data_238 = 8'h0c; // @[Expression.scala 2342:18]
  assign win_data_239 = 8'h0b; // @[Expression.scala 2342:18]
  assign win_data_240 = 8'h0a; // @[Expression.scala 2342:18]
  assign win_data_241 = 8'h09; // @[Expression.scala 2342:18]
  assign win_data_242 = 8'h07; // @[Expression.scala 2342:18]
  assign win_data_243 = 8'h06; // @[Expression.scala 2342:18]
  assign win_data_244 = 8'h05; // @[Expression.scala 2342:18]
  assign win_data_245 = 8'h05; // @[Expression.scala 2342:18]
  assign win_data_246 = 8'h04; // @[Expression.scala 2342:18]
  assign win_data_247 = 8'h03; // @[Expression.scala 2342:18]
  assign win_data_248 = 8'h02; // @[Expression.scala 2342:18]
  assign win_data_249 = 8'h02; // @[Expression.scala 2342:18]
  assign win_data_250 = 8'h01; // @[Expression.scala 2342:18]
  assign win_data_251 = 8'h01; // @[Expression.scala 2342:18]
  assign win_data_252 = 8'h01; // @[Expression.scala 2342:18]
  assign win_data_253 = 8'h0; // @[Expression.scala 2342:18]
  assign win_data_254 = 8'h0; // @[Expression.scala 2342:18]
  assign win_data_255 = 8'h0; // @[Expression.scala 2342:18]
  assign win = tmp_win; // @[win_rom.scala 26:10]

endmodule
